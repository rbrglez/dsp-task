--------------------------------------------------------------------------------
-- fix_matrix_vector_product
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Libraries
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

library olo;
use olo.olo_base_pkg_array.all;
use olo.en_cl_fix_pkg.all;
use olo.olo_fix_pkg.all;

library work;
use work.extend_pkg_array.all;

--------------------------------------------------------------------------------
-- Entity
--------------------------------------------------------------------------------
entity fix_matrix_vector_product is
    generic (
        NUM_DOT_PRODUCTS_G : positive := 11;

        MATRIX_ROW_WIDTH_G    : natural := 32;
        MATRIX_COLUMN_WIDTH_G : natural := 32;

        FMT_IN_MATRIX_ELEMENT_G : string := "(0, 8, 8)";
        FMT_IN_VECTOR_ELEMENT_G : string := "(0, 8, 8)";
        FMT_OUT_RESULT_G        : string := "(0, 21, 16)"
    );
    port (
        clk_i : in std_logic;
        rst_i : in std_logic;

        ------------------------------------------------------------------------
        -- In Interface
        ------------------------------------------------------------------------
        in_valid_i  : in  std_logic := '1';
        in_ready_o  : out std_logic;
        in_matrix_i : in  StlvVectorArray_t(MATRIX_ROW_WIDTH_G - 1 downto 0)(MATRIX_COLUMN_WIDTH_G - 1 downto 0)(fixFmtWidthFromString(FMT_IN_MATRIX_ELEMENT_G) - 1 downto 0);
        in_vector_i : in  StlvArray_t(MATRIX_COLUMN_WIDTH_G - 1 downto 0)(fixFmtWidthFromString(FMT_IN_VECTOR_ELEMENT_G) - 1 downto 0);

        ------------------------------------------------------------------------
        -- Out Interface
        ------------------------------------------------------------------------
        out_valid_o  : out std_logic;
        out_error_o  : out std_logic;
        out_result_o : out StlvArray_t(MATRIX_ROW_WIDTH_G - 1 downto 0)(fixFmtWidthFromString(FMT_OUT_RESULT_G) - 1 downto 0)
    );
end entity fix_matrix_vector_product;

architecture rtl of fix_matrix_vector_product is

    ----------------------------------------------------------------------------
    -- Constants
    ----------------------------------------------------------------------------
    -- Number of fix_dot_product stages needed to compute the final out_result.
    constant NUM_STAGES_C : positive := integer(ceil(real(MATRIX_ROW_WIDTH_G) / real(NUM_DOT_PRODUCTS_G)));

    ----------------------------------------------------------------------------
    -- Types
    ----------------------------------------------------------------------------
    type state_t is (
            IDLE_S,
            FEED_DOT_PRODUCT_S,
            COLLECT_DOT_PRODUCT_S
        );

    type two_process_r is record
        in_ready        : std_logic;
        out_valid       : std_logic;
        out_error       : std_logic;
        out_result      : StlvArray_t(MATRIX_ROW_WIDTH_G - 1 downto 0)(fixFmtWidthFromString(FMT_OUT_RESULT_G) - 1 downto 0);
        in_dot_valid    : std_logic;
        matrix_extended : StlvVectorArray_t(NUM_DOT_PRODUCTS_G*NUM_STAGES_C - 1 downto 0)(MATRIX_COLUMN_WIDTH_G - 1 downto 0)(fixFmtWidthFromString(FMT_IN_MATRIX_ELEMENT_G) - 1 downto 0);
        vector          : StlvArray_t(MATRIX_COLUMN_WIDTH_G - 1 downto 0)(fixFmtWidthFromString(FMT_IN_VECTOR_ELEMENT_G) - 1 downto 0);
        stage_idx       : natural range 0 to NUM_STAGES_C;
        --
        state : state_t;
    end record;

    ----------------------------------------------------------------------------
    -- Two Process records
    ----------------------------------------------------------------------------
    signal r      : two_process_r;
    signal r_next : two_process_r;

    ----------------------------------------------------------------------------
    -- Fix Dot Product signals
    ----------------------------------------------------------------------------
    signal in_dot_ready : std_logic_vector(NUM_DOT_PRODUCTS_G - 1 downto 0);

    signal out_dot_valid  : std_logic_vector(NUM_DOT_PRODUCTS_G - 1 downto 0);
    signal out_dot_result : StlvArray_t(NUM_DOT_PRODUCTS_G - 1 downto 0)(fixFmtWidthFromString(FMT_OUT_RESULT_G) - 1 downto 0);

begin

    ----------------------------------------------------------------------------
    -- Dot Product
    ----------------------------------------------------------------------------
    GEN_DOT_PRODUCT : for i in 0 to NUM_DOT_PRODUCTS_G - 1 generate
        u_fix_dot_product : entity work.fix_dot_product
            generic map (
                DIMENSION_WIDTH_G => MATRIX_COLUMN_WIDTH_G,

                FMT_IN_ELEMENT_A_G => FMT_IN_MATRIX_ELEMENT_G,
                FMT_IN_ELEMENT_B_G => FMT_IN_VECTOR_ELEMENT_G,
                FMT_OUT_RESULT_G   => FMT_OUT_RESULT_G
            )
            port map (
                clk_i => clk_i,
                rst_i => rst_i,

                in_valid_i    => r.in_dot_valid,
                in_ready_o    => in_dot_ready(i),
                in_vector_a_i => r.matrix_extended(i + r.stage_idx * NUM_DOT_PRODUCTS_G),
                in_vector_b_i => r.vector,

                out_valid_o  => out_dot_valid(i),
                out_result_o => out_dot_result(i)
            );
    end generate GEN_DOT_PRODUCT;

    ----------------------------------------------------------------------------
    -- Combinatorial process
    ----------------------------------------------------------------------------
    p_comb : process(all) is
        variable v : two_process_r;
    begin

        -- Hold variables stable
        v := r;

        -- Single clock cycle pulse
        v.out_valid := '0';
        v.out_error := '0';

        ------------------------------------------------------------------------
        -- FSM
        ------------------------------------------------------------------------
        case (r.state) is
            --------------------------------------------------------------------
            when IDLE_S =>
                v.stage_idx := 0;

                v.in_ready := '1';
                if in_valid_i = '1' and r.in_ready = '1' then
                    v.in_ready := '0';

                    -- Register Vector and Matrix
                    v.matrix_extended(MATRIX_ROW_WIDTH_G - 1 downto 0) := in_matrix_i;
                    v.vector                                           := in_vector_i;

                    v.in_dot_valid := '1';
                    v.state        := FEED_DOT_PRODUCT_S;
                end if;

            --------------------------------------------------------------------
            when FEED_DOT_PRODUCT_S =>
                v.in_dot_valid := '1';
                -- Check if in_dot_valid is set and at least one of the
                -- NUM_DOT_PRODUCTS_G fix_dot_product units is ready.
                if (r.in_dot_valid = '1' and in_dot_ready /= (in_dot_ready'range => '0')) then
                    v.in_dot_valid := '0';

                    if (in_dot_ready /= (in_dot_ready'range => '1')) then
                        -- ERROR: 
                        -- All fix_dot_product units must be ready when in_dot_valid is set.
                        v.out_error := '1';
                        v.state     := IDLE_S;
                    else
                        -- Wait for fix_dot_product units to finish computing the dot products.
                        v.state := COLLECT_DOT_PRODUCT_S;
                    end if;
                end if;

            --------------------------------------------------------------------
            when COLLECT_DOT_PRODUCT_S =>

                -- Check if at least one of the NUM_DOT_PRODUCTS_G
                -- fix_dot_product units has out_dot_valid set.
                if (out_dot_valid /= (out_dot_valid'range => '0')) then

                    -- In this stage, populate up to NUM_DOT_PRODUCTS_G elements
                    -- of the result vector with computed dot_product results.
                    for i in 0 to NUM_DOT_PRODUCTS_G - 1 loop
                        if (i + r.stage_idx * NUM_DOT_PRODUCTS_G < MATRIX_ROW_WIDTH_G) then
                            v.out_result(i + r.stage_idx * NUM_DOT_PRODUCTS_G) := out_dot_result(i);
                        end if;
                    end loop;

                    if (out_dot_valid /= (out_dot_valid'range => '1')) then
                        -- ERROR: 
                        -- All fix_dot_product units must set out_dot_valid simultaneously.
                        v.out_error := '1';
                        v.state     := IDLE_S;

                    elsif (r.stage_idx < NUM_STAGES_C - 1) then
                        -- Start a new stage of dot_product calculation
                        v.stage_idx    := r.stage_idx + 1;
                        v.in_dot_valid := '1';
                        v.state        := FEED_DOT_PRODUCT_S;

                    else
                        -- All stages (NUM_STAGES_C) of the dot_product calculation are done. 
                        -- out_result vector contains the complete result.
                        v.out_valid := '1';
                        v.in_ready  := '1';
                        v.stage_idx := 0;
                        v.state     := IDLE_S;
                    end if;
                end if;

            --------------------------------------------------------------------
            when others =>
                null;
        ------------------------------------------------------------------------
        end case;

        -- Apply to record
        r_next <= v;

    end process;

    ----------------------------------------------------------------------------
    -- Output
    ----------------------------------------------------------------------------
    -- In Interface
    in_ready_o <= r.in_ready;
    -- Out Interface
    out_valid_o  <= r.out_valid;
    out_error_o  <= r.out_error;
    out_result_o <= r.out_result;

    ----------------------------------------------------------------------------
    -- Sequential Process
    ----------------------------------------------------------------------------
    p_seq : process(clk_i) is
    begin
        if rising_edge(clk_i) then
            r <= r_next;
            if (rst_i = '1') then
                r.in_ready        <= '1';
                r.out_valid       <= '0';
                r.out_error       <= '0';
                r.in_dot_valid    <= '0';
                r.stage_idx       <= 0;
                r.matrix_extended <= (others => (others => (others => 'X')));
                r.state           <= IDLE_S;
            end if;
        end if;
    end process;

end architecture rtl;
